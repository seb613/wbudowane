-- LAB01SYSWBUDOWANE.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity LAB01SYSWBUDOWANE is
	port (
		clk_clk           : in  std_logic                     := '0';             --        clk.clk
		hex_export        : out std_logic_vector(47 downto 0);                    --        hex.export
		leds_export       : out std_logic_vector(9 downto 0);                     --       leds.export
		pushbutton_export : in  std_logic_vector(3 downto 0)  := (others => '0'); -- pushbutton.export
		reset_reset_n     : in  std_logic                     := '0';             --      reset.reset_n
		sw_sliders_export : in  std_logic_vector(9 downto 0)  := (others => '0')  -- sw_sliders.export
	);
end entity LAB01SYSWBUDOWANE;

architecture rtl of LAB01SYSWBUDOWANE is
	component LAB01SYSWBUDOWANE_HEX is
		port (
			s_address   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			s_read      : in  std_logic                     := 'X';             -- read
			s_readdata  : out std_logic_vector(7 downto 0);                     -- readdata
			s_write     : in  std_logic                     := 'X';             -- write
			s_writedata : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			SEG7        : out std_logic_vector(47 downto 0);                    -- export
			s_clk       : in  std_logic                     := 'X';             -- clk
			s_reset     : in  std_logic                     := 'X'              -- reset
		);
	end component LAB01SYSWBUDOWANE_HEX;

	component LAB01SYSWBUDOWANE_JTAG_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component LAB01SYSWBUDOWANE_JTAG_UART;

	component LAB01SYSWBUDOWANE_NIOS_II_Processor is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(18 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(18 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component LAB01SYSWBUDOWANE_NIOS_II_Processor;

	component LAB01SYSWBUDOWANE_OnChip_Memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component LAB01SYSWBUDOWANE_OnChip_Memory;

	component LAB01SYSWBUDOWANE_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component LAB01SYSWBUDOWANE_leds;

	component LAB01SYSWBUDOWANE_pushbutton is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component LAB01SYSWBUDOWANE_pushbutton;

	component LAB01SYSWBUDOWANE_sw_sliders is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component LAB01SYSWBUDOWANE_sw_sliders;

	component LAB01SYSWBUDOWANE_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                       : in  std_logic                     := 'X';             -- clk
			HEX_clock_sink_reset_reset_bridge_in_reset_reset    : in  std_logic                     := 'X';             -- reset
			NIOS_II_Processor_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			OnChip_Memory_reset1_reset_bridge_in_reset_reset    : in  std_logic                     := 'X';             -- reset
			NIOS_II_Processor_data_master_address               : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			NIOS_II_Processor_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			NIOS_II_Processor_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			NIOS_II_Processor_data_master_read                  : in  std_logic                     := 'X';             -- read
			NIOS_II_Processor_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			NIOS_II_Processor_data_master_readdatavalid         : out std_logic;                                        -- readdatavalid
			NIOS_II_Processor_data_master_write                 : in  std_logic                     := 'X';             -- write
			NIOS_II_Processor_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			NIOS_II_Processor_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			NIOS_II_Processor_instruction_master_address        : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			NIOS_II_Processor_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			NIOS_II_Processor_instruction_master_read           : in  std_logic                     := 'X';             -- read
			NIOS_II_Processor_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			NIOS_II_Processor_instruction_master_readdatavalid  : out std_logic;                                        -- readdatavalid
			HEX_avalon_slave_address                            : out std_logic_vector(2 downto 0);                     -- address
			HEX_avalon_slave_write                              : out std_logic;                                        -- write
			HEX_avalon_slave_read                               : out std_logic;                                        -- read
			HEX_avalon_slave_readdata                           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			HEX_avalon_slave_writedata                          : out std_logic_vector(7 downto 0);                     -- writedata
			JTAG_UART_avalon_jtag_slave_address                 : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_avalon_jtag_slave_write                   : out std_logic;                                        -- write
			JTAG_UART_avalon_jtag_slave_read                    : out std_logic;                                        -- read
			JTAG_UART_avalon_jtag_slave_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_avalon_jtag_slave_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_avalon_jtag_slave_waitrequest             : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect              : out std_logic;                                        -- chipselect
			leds_s1_address                                     : out std_logic_vector(1 downto 0);                     -- address
			leds_s1_write                                       : out std_logic;                                        -- write
			leds_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                                  : out std_logic;                                        -- chipselect
			NIOS_II_Processor_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			NIOS_II_Processor_debug_mem_slave_write             : out std_logic;                                        -- write
			NIOS_II_Processor_debug_mem_slave_read              : out std_logic;                                        -- read
			NIOS_II_Processor_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			NIOS_II_Processor_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			NIOS_II_Processor_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			NIOS_II_Processor_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			NIOS_II_Processor_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			OnChip_Memory_s1_address                            : out std_logic_vector(14 downto 0);                    -- address
			OnChip_Memory_s1_write                              : out std_logic;                                        -- write
			OnChip_Memory_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			OnChip_Memory_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			OnChip_Memory_s1_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			OnChip_Memory_s1_chipselect                         : out std_logic;                                        -- chipselect
			OnChip_Memory_s1_clken                              : out std_logic;                                        -- clken
			pushbutton_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pushbutton_s1_write                                 : out std_logic;                                        -- write
			pushbutton_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pushbutton_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pushbutton_s1_chipselect                            : out std_logic;                                        -- chipselect
			sw_sliders_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			sw_sliders_s1_write                                 : out std_logic;                                        -- write
			sw_sliders_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sw_sliders_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			sw_sliders_s1_chipselect                            : out std_logic                                         -- chipselect
		);
	end component LAB01SYSWBUDOWANE_mm_interconnect_0;

	component LAB01SYSWBUDOWANE_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component LAB01SYSWBUDOWANE_irq_mapper;

	component lab01syswbudowane_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lab01syswbudowane_rst_controller;

	component lab01syswbudowane_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lab01syswbudowane_rst_controller_001;

	component lab01syswbudowane_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lab01syswbudowane_rst_controller_002;

	signal nios_ii_processor_data_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS_II_Processor_data_master_readdata -> NIOS_II_Processor:d_readdata
	signal nios_ii_processor_data_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:NIOS_II_Processor_data_master_waitrequest -> NIOS_II_Processor:d_waitrequest
	signal nios_ii_processor_data_master_debugaccess                       : std_logic;                     -- NIOS_II_Processor:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_II_Processor_data_master_debugaccess
	signal nios_ii_processor_data_master_address                           : std_logic_vector(18 downto 0); -- NIOS_II_Processor:d_address -> mm_interconnect_0:NIOS_II_Processor_data_master_address
	signal nios_ii_processor_data_master_byteenable                        : std_logic_vector(3 downto 0);  -- NIOS_II_Processor:d_byteenable -> mm_interconnect_0:NIOS_II_Processor_data_master_byteenable
	signal nios_ii_processor_data_master_read                              : std_logic;                     -- NIOS_II_Processor:d_read -> mm_interconnect_0:NIOS_II_Processor_data_master_read
	signal nios_ii_processor_data_master_readdatavalid                     : std_logic;                     -- mm_interconnect_0:NIOS_II_Processor_data_master_readdatavalid -> NIOS_II_Processor:d_readdatavalid
	signal nios_ii_processor_data_master_write                             : std_logic;                     -- NIOS_II_Processor:d_write -> mm_interconnect_0:NIOS_II_Processor_data_master_write
	signal nios_ii_processor_data_master_writedata                         : std_logic_vector(31 downto 0); -- NIOS_II_Processor:d_writedata -> mm_interconnect_0:NIOS_II_Processor_data_master_writedata
	signal nios_ii_processor_instruction_master_readdata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS_II_Processor_instruction_master_readdata -> NIOS_II_Processor:i_readdata
	signal nios_ii_processor_instruction_master_waitrequest                : std_logic;                     -- mm_interconnect_0:NIOS_II_Processor_instruction_master_waitrequest -> NIOS_II_Processor:i_waitrequest
	signal nios_ii_processor_instruction_master_address                    : std_logic_vector(18 downto 0); -- NIOS_II_Processor:i_address -> mm_interconnect_0:NIOS_II_Processor_instruction_master_address
	signal nios_ii_processor_instruction_master_read                       : std_logic;                     -- NIOS_II_Processor:i_read -> mm_interconnect_0:NIOS_II_Processor_instruction_master_read
	signal nios_ii_processor_instruction_master_readdatavalid              : std_logic;                     -- mm_interconnect_0:NIOS_II_Processor_instruction_master_readdatavalid -> NIOS_II_Processor:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect        : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata          : std_logic_vector(31 downto 0); -- JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest       : std_logic;                     -- JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address           : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read              : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write             : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	signal mm_interconnect_0_hex_avalon_slave_readdata                     : std_logic_vector(7 downto 0);  -- HEX:s_readdata -> mm_interconnect_0:HEX_avalon_slave_readdata
	signal mm_interconnect_0_hex_avalon_slave_address                      : std_logic_vector(2 downto 0);  -- mm_interconnect_0:HEX_avalon_slave_address -> HEX:s_address
	signal mm_interconnect_0_hex_avalon_slave_read                         : std_logic;                     -- mm_interconnect_0:HEX_avalon_slave_read -> HEX:s_read
	signal mm_interconnect_0_hex_avalon_slave_write                        : std_logic;                     -- mm_interconnect_0:HEX_avalon_slave_write -> HEX:s_write
	signal mm_interconnect_0_hex_avalon_slave_writedata                    : std_logic_vector(7 downto 0);  -- mm_interconnect_0:HEX_avalon_slave_writedata -> HEX:s_writedata
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_readdata    : std_logic_vector(31 downto 0); -- NIOS_II_Processor:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_readdata
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_waitrequest : std_logic;                     -- NIOS_II_Processor:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_debugaccess : std_logic;                     -- mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_debugaccess -> NIOS_II_Processor:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_address     : std_logic_vector(8 downto 0);  -- mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_address -> NIOS_II_Processor:debug_mem_slave_address
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_read        : std_logic;                     -- mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_read -> NIOS_II_Processor:debug_mem_slave_read
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_byteenable -> NIOS_II_Processor:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_write       : std_logic;                     -- mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_write -> NIOS_II_Processor:debug_mem_slave_write
	signal mm_interconnect_0_nios_ii_processor_debug_mem_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_writedata -> NIOS_II_Processor:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:OnChip_Memory_s1_chipselect -> OnChip_Memory:chipselect
	signal mm_interconnect_0_onchip_memory_s1_readdata                     : std_logic_vector(31 downto 0); -- OnChip_Memory:readdata -> mm_interconnect_0:OnChip_Memory_s1_readdata
	signal mm_interconnect_0_onchip_memory_s1_address                      : std_logic_vector(14 downto 0); -- mm_interconnect_0:OnChip_Memory_s1_address -> OnChip_Memory:address
	signal mm_interconnect_0_onchip_memory_s1_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:OnChip_Memory_s1_byteenable -> OnChip_Memory:byteenable
	signal mm_interconnect_0_onchip_memory_s1_write                        : std_logic;                     -- mm_interconnect_0:OnChip_Memory_s1_write -> OnChip_Memory:write
	signal mm_interconnect_0_onchip_memory_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:OnChip_Memory_s1_writedata -> OnChip_Memory:writedata
	signal mm_interconnect_0_onchip_memory_s1_clken                        : std_logic;                     -- mm_interconnect_0:OnChip_Memory_s1_clken -> OnChip_Memory:clken
	signal mm_interconnect_0_leds_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_0_leds_s1_readdata                              : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_0:leds_s1_readdata
	signal mm_interconnect_0_leds_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_s1_address -> leds:address
	signal mm_interconnect_0_leds_s1_write                                 : std_logic;                     -- mm_interconnect_0:leds_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_s1_writedata -> leds:writedata
	signal mm_interconnect_0_sw_sliders_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:sw_sliders_s1_chipselect -> sw_sliders:chipselect
	signal mm_interconnect_0_sw_sliders_s1_readdata                        : std_logic_vector(31 downto 0); -- sw_sliders:readdata -> mm_interconnect_0:sw_sliders_s1_readdata
	signal mm_interconnect_0_sw_sliders_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sw_sliders_s1_address -> sw_sliders:address
	signal mm_interconnect_0_sw_sliders_s1_write                           : std_logic;                     -- mm_interconnect_0:sw_sliders_s1_write -> mm_interconnect_0_sw_sliders_s1_write:in
	signal mm_interconnect_0_sw_sliders_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:sw_sliders_s1_writedata -> sw_sliders:writedata
	signal mm_interconnect_0_pushbutton_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pushbutton_s1_chipselect -> pushbutton:chipselect
	signal mm_interconnect_0_pushbutton_s1_readdata                        : std_logic_vector(31 downto 0); -- pushbutton:readdata -> mm_interconnect_0:pushbutton_s1_readdata
	signal mm_interconnect_0_pushbutton_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pushbutton_s1_address -> pushbutton:address
	signal mm_interconnect_0_pushbutton_s1_write                           : std_logic;                     -- mm_interconnect_0:pushbutton_s1_write -> mm_interconnect_0_pushbutton_s1_write:in
	signal mm_interconnect_0_pushbutton_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pushbutton_s1_writedata -> pushbutton:writedata
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- sw_sliders:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- pushbutton:irq -> irq_mapper:receiver2_irq
	signal nios_ii_processor_irq_irq                                       : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> NIOS_II_Processor:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [HEX:s_reset, mm_interconnect_0:HEX_clock_sink_reset_reset_bridge_in_reset_reset]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:NIOS_II_Processor_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                          : std_logic;                     -- rst_controller_001:reset_req -> [NIOS_II_Processor:reset_req, rst_translator:reset_req_in]
	signal nios_ii_processor_debug_reset_request_reset                     : std_logic;                     -- NIOS_II_Processor:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	signal rst_controller_002_reset_out_reset                              : std_logic;                     -- rst_controller_002:reset_out -> [OnChip_Memory:reset, mm_interconnect_0:OnChip_Memory_reset1_reset_bridge_in_reset_reset]
	signal rst_controller_002_reset_out_reset_req                          : std_logic;                     -- rst_controller_002:reset_req -> OnChip_Memory:reset_req
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv    : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> JTAG_UART:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv   : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> JTAG_UART:av_write_n
	signal mm_interconnect_0_leds_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> leds:write_n
	signal mm_interconnect_0_sw_sliders_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_sw_sliders_s1_write:inv -> sw_sliders:write_n
	signal mm_interconnect_0_pushbutton_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pushbutton_s1_write:inv -> pushbutton:write_n
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [JTAG_UART:rst_n, NIOS_II_Processor:reset_n, leds:reset_n, pushbutton:reset_n, sw_sliders:reset_n]

begin

	hex : component LAB01SYSWBUDOWANE_HEX
		port map (
			s_address   => mm_interconnect_0_hex_avalon_slave_address,   --     avalon_slave.address
			s_read      => mm_interconnect_0_hex_avalon_slave_read,      --                 .read
			s_readdata  => mm_interconnect_0_hex_avalon_slave_readdata,  --                 .readdata
			s_write     => mm_interconnect_0_hex_avalon_slave_write,     --                 .write
			s_writedata => mm_interconnect_0_hex_avalon_slave_writedata, --                 .writedata
			SEG7        => hex_export,                                   --      conduit_end.export
			s_clk       => clk_clk,                                      --       clock_sink.clk
			s_reset     => rst_controller_reset_out_reset                -- clock_sink_reset.reset
		);

	jtag_uart : component LAB01SYSWBUDOWANE_JTAG_UART
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	nios_ii_processor : component LAB01SYSWBUDOWANE_NIOS_II_Processor
		port map (
			clk                                 => clk_clk,                                                         --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,                    --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,                          --                          .reset_req
			d_address                           => nios_ii_processor_data_master_address,                           --               data_master.address
			d_byteenable                        => nios_ii_processor_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios_ii_processor_data_master_read,                              --                          .read
			d_readdata                          => nios_ii_processor_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios_ii_processor_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios_ii_processor_data_master_write,                             --                          .write
			d_writedata                         => nios_ii_processor_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios_ii_processor_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios_ii_processor_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios_ii_processor_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios_ii_processor_instruction_master_read,                       --                          .read
			i_readdata                          => nios_ii_processor_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios_ii_processor_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios_ii_processor_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios_ii_processor_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios_ii_processor_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios_ii_processor_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios_ii_processor_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios_ii_processor_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios_ii_processor_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios_ii_processor_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios_ii_processor_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios_ii_processor_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios_ii_processor_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                             -- custom_instruction_master.readra
		);

	onchip_memory : component LAB01SYSWBUDOWANE_OnChip_Memory
		port map (
			clk        => clk_clk,                                       --   clk1.clk
			address    => mm_interconnect_0_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_002_reset_out_reset,            -- reset1.reset
			reset_req  => rst_controller_002_reset_out_reset_req,        --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	leds : component LAB01SYSWBUDOWANE_leds
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,            --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv,    --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,          --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,         --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,           --                    .readdata
			out_port   => leds_export                                   -- external_connection.export
		);

	pushbutton : component LAB01SYSWBUDOWANE_pushbutton
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_pushbutton_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pushbutton_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pushbutton_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pushbutton_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pushbutton_s1_readdata,        --                    .readdata
			in_port    => pushbutton_export,                               -- external_connection.export
			irq        => irq_mapper_receiver2_irq                         --                 irq.irq
		);

	sw_sliders : component LAB01SYSWBUDOWANE_sw_sliders
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_sw_sliders_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_sw_sliders_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_sw_sliders_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_sw_sliders_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_sw_sliders_s1_readdata,        --                    .readdata
			in_port    => sw_sliders_export,                               -- external_connection.export
			irq        => irq_mapper_receiver1_irq                         --                 irq.irq
		);

	mm_interconnect_0 : component LAB01SYSWBUDOWANE_mm_interconnect_0
		port map (
			clk_0_clk_clk                                       => clk_clk,                                                         --                                     clk_0_clk.clk
			HEX_clock_sink_reset_reset_bridge_in_reset_reset    => rst_controller_reset_out_reset,                                  --    HEX_clock_sink_reset_reset_bridge_in_reset.reset
			NIOS_II_Processor_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                              -- NIOS_II_Processor_reset_reset_bridge_in_reset.reset
			OnChip_Memory_reset1_reset_bridge_in_reset_reset    => rst_controller_002_reset_out_reset,                              --    OnChip_Memory_reset1_reset_bridge_in_reset.reset
			NIOS_II_Processor_data_master_address               => nios_ii_processor_data_master_address,                           --                 NIOS_II_Processor_data_master.address
			NIOS_II_Processor_data_master_waitrequest           => nios_ii_processor_data_master_waitrequest,                       --                                              .waitrequest
			NIOS_II_Processor_data_master_byteenable            => nios_ii_processor_data_master_byteenable,                        --                                              .byteenable
			NIOS_II_Processor_data_master_read                  => nios_ii_processor_data_master_read,                              --                                              .read
			NIOS_II_Processor_data_master_readdata              => nios_ii_processor_data_master_readdata,                          --                                              .readdata
			NIOS_II_Processor_data_master_readdatavalid         => nios_ii_processor_data_master_readdatavalid,                     --                                              .readdatavalid
			NIOS_II_Processor_data_master_write                 => nios_ii_processor_data_master_write,                             --                                              .write
			NIOS_II_Processor_data_master_writedata             => nios_ii_processor_data_master_writedata,                         --                                              .writedata
			NIOS_II_Processor_data_master_debugaccess           => nios_ii_processor_data_master_debugaccess,                       --                                              .debugaccess
			NIOS_II_Processor_instruction_master_address        => nios_ii_processor_instruction_master_address,                    --          NIOS_II_Processor_instruction_master.address
			NIOS_II_Processor_instruction_master_waitrequest    => nios_ii_processor_instruction_master_waitrequest,                --                                              .waitrequest
			NIOS_II_Processor_instruction_master_read           => nios_ii_processor_instruction_master_read,                       --                                              .read
			NIOS_II_Processor_instruction_master_readdata       => nios_ii_processor_instruction_master_readdata,                   --                                              .readdata
			NIOS_II_Processor_instruction_master_readdatavalid  => nios_ii_processor_instruction_master_readdatavalid,              --                                              .readdatavalid
			HEX_avalon_slave_address                            => mm_interconnect_0_hex_avalon_slave_address,                      --                              HEX_avalon_slave.address
			HEX_avalon_slave_write                              => mm_interconnect_0_hex_avalon_slave_write,                        --                                              .write
			HEX_avalon_slave_read                               => mm_interconnect_0_hex_avalon_slave_read,                         --                                              .read
			HEX_avalon_slave_readdata                           => mm_interconnect_0_hex_avalon_slave_readdata,                     --                                              .readdata
			HEX_avalon_slave_writedata                          => mm_interconnect_0_hex_avalon_slave_writedata,                    --                                              .writedata
			JTAG_UART_avalon_jtag_slave_address                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,           --                   JTAG_UART_avalon_jtag_slave.address
			JTAG_UART_avalon_jtag_slave_write                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,             --                                              .write
			JTAG_UART_avalon_jtag_slave_read                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,              --                                              .read
			JTAG_UART_avalon_jtag_slave_readdata                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,          --                                              .readdata
			JTAG_UART_avalon_jtag_slave_writedata               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,         --                                              .writedata
			JTAG_UART_avalon_jtag_slave_waitrequest             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,       --                                              .waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect              => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,        --                                              .chipselect
			leds_s1_address                                     => mm_interconnect_0_leds_s1_address,                               --                                       leds_s1.address
			leds_s1_write                                       => mm_interconnect_0_leds_s1_write,                                 --                                              .write
			leds_s1_readdata                                    => mm_interconnect_0_leds_s1_readdata,                              --                                              .readdata
			leds_s1_writedata                                   => mm_interconnect_0_leds_s1_writedata,                             --                                              .writedata
			leds_s1_chipselect                                  => mm_interconnect_0_leds_s1_chipselect,                            --                                              .chipselect
			NIOS_II_Processor_debug_mem_slave_address           => mm_interconnect_0_nios_ii_processor_debug_mem_slave_address,     --             NIOS_II_Processor_debug_mem_slave.address
			NIOS_II_Processor_debug_mem_slave_write             => mm_interconnect_0_nios_ii_processor_debug_mem_slave_write,       --                                              .write
			NIOS_II_Processor_debug_mem_slave_read              => mm_interconnect_0_nios_ii_processor_debug_mem_slave_read,        --                                              .read
			NIOS_II_Processor_debug_mem_slave_readdata          => mm_interconnect_0_nios_ii_processor_debug_mem_slave_readdata,    --                                              .readdata
			NIOS_II_Processor_debug_mem_slave_writedata         => mm_interconnect_0_nios_ii_processor_debug_mem_slave_writedata,   --                                              .writedata
			NIOS_II_Processor_debug_mem_slave_byteenable        => mm_interconnect_0_nios_ii_processor_debug_mem_slave_byteenable,  --                                              .byteenable
			NIOS_II_Processor_debug_mem_slave_waitrequest       => mm_interconnect_0_nios_ii_processor_debug_mem_slave_waitrequest, --                                              .waitrequest
			NIOS_II_Processor_debug_mem_slave_debugaccess       => mm_interconnect_0_nios_ii_processor_debug_mem_slave_debugaccess, --                                              .debugaccess
			OnChip_Memory_s1_address                            => mm_interconnect_0_onchip_memory_s1_address,                      --                              OnChip_Memory_s1.address
			OnChip_Memory_s1_write                              => mm_interconnect_0_onchip_memory_s1_write,                        --                                              .write
			OnChip_Memory_s1_readdata                           => mm_interconnect_0_onchip_memory_s1_readdata,                     --                                              .readdata
			OnChip_Memory_s1_writedata                          => mm_interconnect_0_onchip_memory_s1_writedata,                    --                                              .writedata
			OnChip_Memory_s1_byteenable                         => mm_interconnect_0_onchip_memory_s1_byteenable,                   --                                              .byteenable
			OnChip_Memory_s1_chipselect                         => mm_interconnect_0_onchip_memory_s1_chipselect,                   --                                              .chipselect
			OnChip_Memory_s1_clken                              => mm_interconnect_0_onchip_memory_s1_clken,                        --                                              .clken
			pushbutton_s1_address                               => mm_interconnect_0_pushbutton_s1_address,                         --                                 pushbutton_s1.address
			pushbutton_s1_write                                 => mm_interconnect_0_pushbutton_s1_write,                           --                                              .write
			pushbutton_s1_readdata                              => mm_interconnect_0_pushbutton_s1_readdata,                        --                                              .readdata
			pushbutton_s1_writedata                             => mm_interconnect_0_pushbutton_s1_writedata,                       --                                              .writedata
			pushbutton_s1_chipselect                            => mm_interconnect_0_pushbutton_s1_chipselect,                      --                                              .chipselect
			sw_sliders_s1_address                               => mm_interconnect_0_sw_sliders_s1_address,                         --                                 sw_sliders_s1.address
			sw_sliders_s1_write                                 => mm_interconnect_0_sw_sliders_s1_write,                           --                                              .write
			sw_sliders_s1_readdata                              => mm_interconnect_0_sw_sliders_s1_readdata,                        --                                              .readdata
			sw_sliders_s1_writedata                             => mm_interconnect_0_sw_sliders_s1_writedata,                       --                                              .writedata
			sw_sliders_s1_chipselect                            => mm_interconnect_0_sw_sliders_s1_chipselect                       --                                              .chipselect
		);

	irq_mapper : component LAB01SYSWBUDOWANE_irq_mapper
		port map (
			clk           => clk_clk,                            --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			sender_irq    => nios_ii_processor_irq_irq           --    sender.irq
		);

	rst_controller : component lab01syswbudowane_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component lab01syswbudowane_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                     -- reset_in0.reset
			reset_in1      => nios_ii_processor_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                     --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,          -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req,      --          .reset_req
			reset_req_in0  => '0',                                         -- (terminated)
			reset_req_in1  => '0',                                         -- (terminated)
			reset_in2      => '0',                                         -- (terminated)
			reset_req_in2  => '0',                                         -- (terminated)
			reset_in3      => '0',                                         -- (terminated)
			reset_req_in3  => '0',                                         -- (terminated)
			reset_in4      => '0',                                         -- (terminated)
			reset_req_in4  => '0',                                         -- (terminated)
			reset_in5      => '0',                                         -- (terminated)
			reset_req_in5  => '0',                                         -- (terminated)
			reset_in6      => '0',                                         -- (terminated)
			reset_req_in6  => '0',                                         -- (terminated)
			reset_in7      => '0',                                         -- (terminated)
			reset_req_in7  => '0',                                         -- (terminated)
			reset_in8      => '0',                                         -- (terminated)
			reset_req_in8  => '0',                                         -- (terminated)
			reset_in9      => '0',                                         -- (terminated)
			reset_req_in9  => '0',                                         -- (terminated)
			reset_in10     => '0',                                         -- (terminated)
			reset_req_in10 => '0',                                         -- (terminated)
			reset_in11     => '0',                                         -- (terminated)
			reset_req_in11 => '0',                                         -- (terminated)
			reset_in12     => '0',                                         -- (terminated)
			reset_req_in12 => '0',                                         -- (terminated)
			reset_in13     => '0',                                         -- (terminated)
			reset_req_in13 => '0',                                         -- (terminated)
			reset_in14     => '0',                                         -- (terminated)
			reset_req_in14 => '0',                                         -- (terminated)
			reset_in15     => '0',                                         -- (terminated)
			reset_req_in15 => '0'                                          -- (terminated)
		);

	rst_controller_002 : component lab01syswbudowane_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios_ii_processor_debug_reset_request_reset, -- reset_in0.reset
			clk            => clk_clk,                                     --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,          -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req,      --          .reset_req
			reset_req_in0  => '0',                                         -- (terminated)
			reset_in1      => '0',                                         -- (terminated)
			reset_req_in1  => '0',                                         -- (terminated)
			reset_in2      => '0',                                         -- (terminated)
			reset_req_in2  => '0',                                         -- (terminated)
			reset_in3      => '0',                                         -- (terminated)
			reset_req_in3  => '0',                                         -- (terminated)
			reset_in4      => '0',                                         -- (terminated)
			reset_req_in4  => '0',                                         -- (terminated)
			reset_in5      => '0',                                         -- (terminated)
			reset_req_in5  => '0',                                         -- (terminated)
			reset_in6      => '0',                                         -- (terminated)
			reset_req_in6  => '0',                                         -- (terminated)
			reset_in7      => '0',                                         -- (terminated)
			reset_req_in7  => '0',                                         -- (terminated)
			reset_in8      => '0',                                         -- (terminated)
			reset_req_in8  => '0',                                         -- (terminated)
			reset_in9      => '0',                                         -- (terminated)
			reset_req_in9  => '0',                                         -- (terminated)
			reset_in10     => '0',                                         -- (terminated)
			reset_req_in10 => '0',                                         -- (terminated)
			reset_in11     => '0',                                         -- (terminated)
			reset_req_in11 => '0',                                         -- (terminated)
			reset_in12     => '0',                                         -- (terminated)
			reset_req_in12 => '0',                                         -- (terminated)
			reset_in13     => '0',                                         -- (terminated)
			reset_req_in13 => '0',                                         -- (terminated)
			reset_in14     => '0',                                         -- (terminated)
			reset_req_in14 => '0',                                         -- (terminated)
			reset_in15     => '0',                                         -- (terminated)
			reset_req_in15 => '0'                                          -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	mm_interconnect_0_sw_sliders_s1_write_ports_inv <= not mm_interconnect_0_sw_sliders_s1_write;

	mm_interconnect_0_pushbutton_s1_write_ports_inv <= not mm_interconnect_0_pushbutton_s1_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of LAB01SYSWBUDOWANE
