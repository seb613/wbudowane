// SyswbLab1.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module SyswbLab1 (
		input  wire        clk_clk,           //        clk.clk
		output wire [47:0] hex_export,        //        hex.export
		output wire [9:0]  leds_export,       //       leds.export
		input  wire [3:0]  pushbutton_export, // pushbutton.export
		input  wire        reset_reset_n,     //      reset.reset_n
		input  wire [9:0]  sw_sliders_export  // sw_sliders.export
	);

	wire  [31:0] nios_ii_processor_data_master_readdata;                          // mm_interconnect_0:NIOS_II_Processor_data_master_readdata -> NIOS_II_Processor:d_readdata
	wire         nios_ii_processor_data_master_waitrequest;                       // mm_interconnect_0:NIOS_II_Processor_data_master_waitrequest -> NIOS_II_Processor:d_waitrequest
	wire         nios_ii_processor_data_master_debugaccess;                       // NIOS_II_Processor:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_II_Processor_data_master_debugaccess
	wire  [18:0] nios_ii_processor_data_master_address;                           // NIOS_II_Processor:d_address -> mm_interconnect_0:NIOS_II_Processor_data_master_address
	wire   [3:0] nios_ii_processor_data_master_byteenable;                        // NIOS_II_Processor:d_byteenable -> mm_interconnect_0:NIOS_II_Processor_data_master_byteenable
	wire         nios_ii_processor_data_master_read;                              // NIOS_II_Processor:d_read -> mm_interconnect_0:NIOS_II_Processor_data_master_read
	wire         nios_ii_processor_data_master_write;                             // NIOS_II_Processor:d_write -> mm_interconnect_0:NIOS_II_Processor_data_master_write
	wire  [31:0] nios_ii_processor_data_master_writedata;                         // NIOS_II_Processor:d_writedata -> mm_interconnect_0:NIOS_II_Processor_data_master_writedata
	wire  [31:0] nios_ii_processor_instruction_master_readdata;                   // mm_interconnect_0:NIOS_II_Processor_instruction_master_readdata -> NIOS_II_Processor:i_readdata
	wire         nios_ii_processor_instruction_master_waitrequest;                // mm_interconnect_0:NIOS_II_Processor_instruction_master_waitrequest -> NIOS_II_Processor:i_waitrequest
	wire  [18:0] nios_ii_processor_instruction_master_address;                    // NIOS_II_Processor:i_address -> mm_interconnect_0:NIOS_II_Processor_instruction_master_address
	wire         nios_ii_processor_instruction_master_read;                       // NIOS_II_Processor:i_read -> mm_interconnect_0:NIOS_II_Processor_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;        // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;          // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;       // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;           // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;              // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;             // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;         // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire   [7:0] mm_interconnect_0_hex_avalon_slave_readdata;                     // HEX:s_readdata -> mm_interconnect_0:HEX_avalon_slave_readdata
	wire   [2:0] mm_interconnect_0_hex_avalon_slave_address;                      // mm_interconnect_0:HEX_avalon_slave_address -> HEX:s_address
	wire         mm_interconnect_0_hex_avalon_slave_read;                         // mm_interconnect_0:HEX_avalon_slave_read -> HEX:s_read
	wire         mm_interconnect_0_hex_avalon_slave_write;                        // mm_interconnect_0:HEX_avalon_slave_write -> HEX:s_write
	wire   [7:0] mm_interconnect_0_hex_avalon_slave_writedata;                    // mm_interconnect_0:HEX_avalon_slave_writedata -> HEX:s_writedata
	wire  [31:0] mm_interconnect_0_nios_ii_processor_debug_mem_slave_readdata;    // NIOS_II_Processor:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_ii_processor_debug_mem_slave_waitrequest; // NIOS_II_Processor:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_ii_processor_debug_mem_slave_debugaccess; // mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_debugaccess -> NIOS_II_Processor:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_ii_processor_debug_mem_slave_address;     // mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_address -> NIOS_II_Processor:debug_mem_slave_address
	wire         mm_interconnect_0_nios_ii_processor_debug_mem_slave_read;        // mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_read -> NIOS_II_Processor:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_ii_processor_debug_mem_slave_byteenable;  // mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_byteenable -> NIOS_II_Processor:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_ii_processor_debug_mem_slave_write;       // mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_write -> NIOS_II_Processor:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_ii_processor_debug_mem_slave_writedata;   // mm_interconnect_0:NIOS_II_Processor_debug_mem_slave_writedata -> NIOS_II_Processor:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                   // mm_interconnect_0:OnChip_Memory_s1_chipselect -> OnChip_Memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                     // OnChip_Memory:readdata -> mm_interconnect_0:OnChip_Memory_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory_s1_address;                      // mm_interconnect_0:OnChip_Memory_s1_address -> OnChip_Memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                   // mm_interconnect_0:OnChip_Memory_s1_byteenable -> OnChip_Memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                        // mm_interconnect_0:OnChip_Memory_s1_write -> OnChip_Memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                    // mm_interconnect_0:OnChip_Memory_s1_writedata -> OnChip_Memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                        // mm_interconnect_0:OnChip_Memory_s1_clken -> OnChip_Memory:clken
	wire         mm_interconnect_0_leds_s1_chipselect;                            // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                              // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                               // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                                 // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                             // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_sw_sliders_s1_chipselect;                      // mm_interconnect_0:sw_sliders_s1_chipselect -> sw_sliders:chipselect
	wire  [31:0] mm_interconnect_0_sw_sliders_s1_readdata;                        // sw_sliders:readdata -> mm_interconnect_0:sw_sliders_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_sliders_s1_address;                         // mm_interconnect_0:sw_sliders_s1_address -> sw_sliders:address
	wire         mm_interconnect_0_sw_sliders_s1_write;                           // mm_interconnect_0:sw_sliders_s1_write -> sw_sliders:write_n
	wire  [31:0] mm_interconnect_0_sw_sliders_s1_writedata;                       // mm_interconnect_0:sw_sliders_s1_writedata -> sw_sliders:writedata
	wire         mm_interconnect_0_pushbutton_s1_chipselect;                      // mm_interconnect_0:pushbutton_s1_chipselect -> pushbutton:chipselect
	wire  [31:0] mm_interconnect_0_pushbutton_s1_readdata;                        // pushbutton:readdata -> mm_interconnect_0:pushbutton_s1_readdata
	wire   [1:0] mm_interconnect_0_pushbutton_s1_address;                         // mm_interconnect_0:pushbutton_s1_address -> pushbutton:address
	wire         mm_interconnect_0_pushbutton_s1_write;                           // mm_interconnect_0:pushbutton_s1_write -> pushbutton:write_n
	wire  [31:0] mm_interconnect_0_pushbutton_s1_writedata;                       // mm_interconnect_0:pushbutton_s1_writedata -> pushbutton:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                         // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                           // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                            // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                              // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                          // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         irq_mapper_receiver0_irq;                                        // JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                        // pushbutton:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                        // sw_sliders:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                        // timer_0:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios_ii_processor_irq_irq;                                       // irq_mapper:sender_irq -> NIOS_II_Processor:irq
	wire         rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [HEX:s_reset, mm_interconnect_0:HEX_clock_sink_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                              // rst_controller_001:reset_out -> [JTAG_UART:rst_n, NIOS_II_Processor:reset_n, irq_mapper:reset, leds:reset_n, mm_interconnect_0:NIOS_II_Processor_reset_reset_bridge_in_reset_reset, pushbutton:reset_n, rst_translator:in_reset, sw_sliders:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                          // rst_controller_001:reset_req -> [NIOS_II_Processor:reset_req, rst_translator:reset_req_in]
	wire         nios_ii_processor_debug_reset_request_reset;                     // NIOS_II_Processor:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	wire         rst_controller_002_reset_out_reset;                              // rst_controller_002:reset_out -> [OnChip_Memory:reset, mm_interconnect_0:OnChip_Memory_reset1_reset_bridge_in_reset_reset, timer_0:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                          // rst_controller_002:reset_req -> [OnChip_Memory:reset_req, rst_translator_001:reset_req_in]

	SEG7_IF #(
		.SEG7_NUM       (6),
		.ADDR_WIDTH     (3),
		.DEFAULT_ACTIVE (1),
		.LOW_ACTIVE     (1)
	) hex (
		.s_address   (mm_interconnect_0_hex_avalon_slave_address),   //     avalon_slave.address
		.s_read      (mm_interconnect_0_hex_avalon_slave_read),      //                 .read
		.s_readdata  (mm_interconnect_0_hex_avalon_slave_readdata),  //                 .readdata
		.s_write     (mm_interconnect_0_hex_avalon_slave_write),     //                 .write
		.s_writedata (mm_interconnect_0_hex_avalon_slave_writedata), //                 .writedata
		.SEG7        (hex_export),                                   //      conduit_end.export
		.s_clk       (clk_clk),                                      //       clock_sink.clk
		.s_reset     (rst_controller_reset_out_reset)                // clock_sink_reset.reset
	);

	SyswbLab1_JTAG_UART jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	SyswbLab1_NIOS_II_Processor nios_ii_processor (
		.clk                                 (clk_clk),                                                         //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                             //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                          //                          .reset_req
		.d_address                           (nios_ii_processor_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_ii_processor_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_ii_processor_data_master_read),                              //                          .read
		.d_readdata                          (nios_ii_processor_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_ii_processor_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_ii_processor_data_master_write),                             //                          .write
		.d_writedata                         (nios_ii_processor_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_ii_processor_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_ii_processor_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_ii_processor_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_ii_processor_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_ii_processor_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_ii_processor_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_ii_processor_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_ii_processor_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_ii_processor_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_ii_processor_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_ii_processor_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_ii_processor_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_ii_processor_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_ii_processor_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_ii_processor_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                                 // custom_instruction_master.readra
	);

	SyswbLab1_OnChip_Memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req),        //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	SyswbLab1_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	SyswbLab1_pushbutton pushbutton (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pushbutton_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pushbutton_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pushbutton_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pushbutton_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pushbutton_s1_readdata),   //                    .readdata
		.in_port    (pushbutton_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                    //                 irq.irq
	);

	SyswbLab1_sw_sliders sw_sliders (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_sw_sliders_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sw_sliders_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sw_sliders_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sw_sliders_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sw_sliders_s1_readdata),   //                    .readdata
		.in_port    (sw_sliders_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                    //                 irq.irq
	);

	SyswbLab1_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	SyswbLab1_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                       (clk_clk),                                                         //                                     clk_0_clk.clk
		.HEX_clock_sink_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                                  //    HEX_clock_sink_reset_reset_bridge_in_reset.reset
		.NIOS_II_Processor_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                              // NIOS_II_Processor_reset_reset_bridge_in_reset.reset
		.OnChip_Memory_reset1_reset_bridge_in_reset_reset    (rst_controller_002_reset_out_reset),                              //    OnChip_Memory_reset1_reset_bridge_in_reset.reset
		.NIOS_II_Processor_data_master_address               (nios_ii_processor_data_master_address),                           //                 NIOS_II_Processor_data_master.address
		.NIOS_II_Processor_data_master_waitrequest           (nios_ii_processor_data_master_waitrequest),                       //                                              .waitrequest
		.NIOS_II_Processor_data_master_byteenable            (nios_ii_processor_data_master_byteenable),                        //                                              .byteenable
		.NIOS_II_Processor_data_master_read                  (nios_ii_processor_data_master_read),                              //                                              .read
		.NIOS_II_Processor_data_master_readdata              (nios_ii_processor_data_master_readdata),                          //                                              .readdata
		.NIOS_II_Processor_data_master_write                 (nios_ii_processor_data_master_write),                             //                                              .write
		.NIOS_II_Processor_data_master_writedata             (nios_ii_processor_data_master_writedata),                         //                                              .writedata
		.NIOS_II_Processor_data_master_debugaccess           (nios_ii_processor_data_master_debugaccess),                       //                                              .debugaccess
		.NIOS_II_Processor_instruction_master_address        (nios_ii_processor_instruction_master_address),                    //          NIOS_II_Processor_instruction_master.address
		.NIOS_II_Processor_instruction_master_waitrequest    (nios_ii_processor_instruction_master_waitrequest),                //                                              .waitrequest
		.NIOS_II_Processor_instruction_master_read           (nios_ii_processor_instruction_master_read),                       //                                              .read
		.NIOS_II_Processor_instruction_master_readdata       (nios_ii_processor_instruction_master_readdata),                   //                                              .readdata
		.HEX_avalon_slave_address                            (mm_interconnect_0_hex_avalon_slave_address),                      //                              HEX_avalon_slave.address
		.HEX_avalon_slave_write                              (mm_interconnect_0_hex_avalon_slave_write),                        //                                              .write
		.HEX_avalon_slave_read                               (mm_interconnect_0_hex_avalon_slave_read),                         //                                              .read
		.HEX_avalon_slave_readdata                           (mm_interconnect_0_hex_avalon_slave_readdata),                     //                                              .readdata
		.HEX_avalon_slave_writedata                          (mm_interconnect_0_hex_avalon_slave_writedata),                    //                                              .writedata
		.JTAG_UART_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),           //                   JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),             //                                              .write
		.JTAG_UART_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),              //                                              .read
		.JTAG_UART_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),          //                                              .readdata
		.JTAG_UART_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),         //                                              .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),       //                                              .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),        //                                              .chipselect
		.leds_s1_address                                     (mm_interconnect_0_leds_s1_address),                               //                                       leds_s1.address
		.leds_s1_write                                       (mm_interconnect_0_leds_s1_write),                                 //                                              .write
		.leds_s1_readdata                                    (mm_interconnect_0_leds_s1_readdata),                              //                                              .readdata
		.leds_s1_writedata                                   (mm_interconnect_0_leds_s1_writedata),                             //                                              .writedata
		.leds_s1_chipselect                                  (mm_interconnect_0_leds_s1_chipselect),                            //                                              .chipselect
		.NIOS_II_Processor_debug_mem_slave_address           (mm_interconnect_0_nios_ii_processor_debug_mem_slave_address),     //             NIOS_II_Processor_debug_mem_slave.address
		.NIOS_II_Processor_debug_mem_slave_write             (mm_interconnect_0_nios_ii_processor_debug_mem_slave_write),       //                                              .write
		.NIOS_II_Processor_debug_mem_slave_read              (mm_interconnect_0_nios_ii_processor_debug_mem_slave_read),        //                                              .read
		.NIOS_II_Processor_debug_mem_slave_readdata          (mm_interconnect_0_nios_ii_processor_debug_mem_slave_readdata),    //                                              .readdata
		.NIOS_II_Processor_debug_mem_slave_writedata         (mm_interconnect_0_nios_ii_processor_debug_mem_slave_writedata),   //                                              .writedata
		.NIOS_II_Processor_debug_mem_slave_byteenable        (mm_interconnect_0_nios_ii_processor_debug_mem_slave_byteenable),  //                                              .byteenable
		.NIOS_II_Processor_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_ii_processor_debug_mem_slave_waitrequest), //                                              .waitrequest
		.NIOS_II_Processor_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_ii_processor_debug_mem_slave_debugaccess), //                                              .debugaccess
		.OnChip_Memory_s1_address                            (mm_interconnect_0_onchip_memory_s1_address),                      //                              OnChip_Memory_s1.address
		.OnChip_Memory_s1_write                              (mm_interconnect_0_onchip_memory_s1_write),                        //                                              .write
		.OnChip_Memory_s1_readdata                           (mm_interconnect_0_onchip_memory_s1_readdata),                     //                                              .readdata
		.OnChip_Memory_s1_writedata                          (mm_interconnect_0_onchip_memory_s1_writedata),                    //                                              .writedata
		.OnChip_Memory_s1_byteenable                         (mm_interconnect_0_onchip_memory_s1_byteenable),                   //                                              .byteenable
		.OnChip_Memory_s1_chipselect                         (mm_interconnect_0_onchip_memory_s1_chipselect),                   //                                              .chipselect
		.OnChip_Memory_s1_clken                              (mm_interconnect_0_onchip_memory_s1_clken),                        //                                              .clken
		.pushbutton_s1_address                               (mm_interconnect_0_pushbutton_s1_address),                         //                                 pushbutton_s1.address
		.pushbutton_s1_write                                 (mm_interconnect_0_pushbutton_s1_write),                           //                                              .write
		.pushbutton_s1_readdata                              (mm_interconnect_0_pushbutton_s1_readdata),                        //                                              .readdata
		.pushbutton_s1_writedata                             (mm_interconnect_0_pushbutton_s1_writedata),                       //                                              .writedata
		.pushbutton_s1_chipselect                            (mm_interconnect_0_pushbutton_s1_chipselect),                      //                                              .chipselect
		.sw_sliders_s1_address                               (mm_interconnect_0_sw_sliders_s1_address),                         //                                 sw_sliders_s1.address
		.sw_sliders_s1_write                                 (mm_interconnect_0_sw_sliders_s1_write),                           //                                              .write
		.sw_sliders_s1_readdata                              (mm_interconnect_0_sw_sliders_s1_readdata),                        //                                              .readdata
		.sw_sliders_s1_writedata                             (mm_interconnect_0_sw_sliders_s1_writedata),                       //                                              .writedata
		.sw_sliders_s1_chipselect                            (mm_interconnect_0_sw_sliders_s1_chipselect),                      //                                              .chipselect
		.timer_0_s1_address                                  (mm_interconnect_0_timer_0_s1_address),                            //                                    timer_0_s1.address
		.timer_0_s1_write                                    (mm_interconnect_0_timer_0_s1_write),                              //                                              .write
		.timer_0_s1_readdata                                 (mm_interconnect_0_timer_0_s1_readdata),                           //                                              .readdata
		.timer_0_s1_writedata                                (mm_interconnect_0_timer_0_s1_writedata),                          //                                              .writedata
		.timer_0_s1_chipselect                               (mm_interconnect_0_timer_0_s1_chipselect)                          //                                              .chipselect
	);

	SyswbLab1_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios_ii_processor_irq_irq)           //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                              // reset_in0.reset
		.reset_in1      (nios_ii_processor_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                     //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),          // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req),      //          .reset_req
		.reset_req_in0  (1'b0),                                        // (terminated)
		.reset_req_in1  (1'b0),                                        // (terminated)
		.reset_in2      (1'b0),                                        // (terminated)
		.reset_req_in2  (1'b0),                                        // (terminated)
		.reset_in3      (1'b0),                                        // (terminated)
		.reset_req_in3  (1'b0),                                        // (terminated)
		.reset_in4      (1'b0),                                        // (terminated)
		.reset_req_in4  (1'b0),                                        // (terminated)
		.reset_in5      (1'b0),                                        // (terminated)
		.reset_req_in5  (1'b0),                                        // (terminated)
		.reset_in6      (1'b0),                                        // (terminated)
		.reset_req_in6  (1'b0),                                        // (terminated)
		.reset_in7      (1'b0),                                        // (terminated)
		.reset_req_in7  (1'b0),                                        // (terminated)
		.reset_in8      (1'b0),                                        // (terminated)
		.reset_req_in8  (1'b0),                                        // (terminated)
		.reset_in9      (1'b0),                                        // (terminated)
		.reset_req_in9  (1'b0),                                        // (terminated)
		.reset_in10     (1'b0),                                        // (terminated)
		.reset_req_in10 (1'b0),                                        // (terminated)
		.reset_in11     (1'b0),                                        // (terminated)
		.reset_req_in11 (1'b0),                                        // (terminated)
		.reset_in12     (1'b0),                                        // (terminated)
		.reset_req_in12 (1'b0),                                        // (terminated)
		.reset_in13     (1'b0),                                        // (terminated)
		.reset_req_in13 (1'b0),                                        // (terminated)
		.reset_in14     (1'b0),                                        // (terminated)
		.reset_req_in14 (1'b0),                                        // (terminated)
		.reset_in15     (1'b0),                                        // (terminated)
		.reset_req_in15 (1'b0)                                         // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (nios_ii_processor_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                     //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),          // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req),      //          .reset_req
		.reset_req_in0  (1'b0),                                        // (terminated)
		.reset_in1      (1'b0),                                        // (terminated)
		.reset_req_in1  (1'b0),                                        // (terminated)
		.reset_in2      (1'b0),                                        // (terminated)
		.reset_req_in2  (1'b0),                                        // (terminated)
		.reset_in3      (1'b0),                                        // (terminated)
		.reset_req_in3  (1'b0),                                        // (terminated)
		.reset_in4      (1'b0),                                        // (terminated)
		.reset_req_in4  (1'b0),                                        // (terminated)
		.reset_in5      (1'b0),                                        // (terminated)
		.reset_req_in5  (1'b0),                                        // (terminated)
		.reset_in6      (1'b0),                                        // (terminated)
		.reset_req_in6  (1'b0),                                        // (terminated)
		.reset_in7      (1'b0),                                        // (terminated)
		.reset_req_in7  (1'b0),                                        // (terminated)
		.reset_in8      (1'b0),                                        // (terminated)
		.reset_req_in8  (1'b0),                                        // (terminated)
		.reset_in9      (1'b0),                                        // (terminated)
		.reset_req_in9  (1'b0),                                        // (terminated)
		.reset_in10     (1'b0),                                        // (terminated)
		.reset_req_in10 (1'b0),                                        // (terminated)
		.reset_in11     (1'b0),                                        // (terminated)
		.reset_req_in11 (1'b0),                                        // (terminated)
		.reset_in12     (1'b0),                                        // (terminated)
		.reset_req_in12 (1'b0),                                        // (terminated)
		.reset_in13     (1'b0),                                        // (terminated)
		.reset_req_in13 (1'b0),                                        // (terminated)
		.reset_in14     (1'b0),                                        // (terminated)
		.reset_req_in14 (1'b0),                                        // (terminated)
		.reset_in15     (1'b0),                                        // (terminated)
		.reset_req_in15 (1'b0)                                         // (terminated)
	);

endmodule
